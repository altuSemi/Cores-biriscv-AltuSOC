`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/core/biriscv_defs.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/core/biriscv_decode.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/core/biriscv_decoder.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/core/biriscv_csr.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/core/biriscv_csr_regfile.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/core/biriscv_alu.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/core/biriscv_npc.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/core/biriscv_multiplier.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/core/biriscv_mmu.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/core/biriscv_lsu.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/core/biriscv_issue.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/core/biriscv_frontend.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/core/biriscv_fetch.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/core/biriscv_exec.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/core/biriscv_divider.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/core/riscv_core.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/core/biriscv_xilinx_2r1w.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/core/biriscv_trace_sim.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/core/biriscv_regfile.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/core/biriscv_pipe_ctrl.v"

`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/icache/icache.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/icache/icache_tag_ram.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/icache/icache_data_ram.v"

`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/dcache/dcache.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/dcache/dcache_axi.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/dcache/dcache_pmem_mux.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/dcache/dcache_mux.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/dcache/dcache_if_pmem.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/dcache/dcache_core.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/dcache/dcache_core_tag_ram.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/dcache/dcache_core_tag_ram.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/dcache/dcache_core_data_ram.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/dcache/dcache_axi_axi.v"

`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/top/riscv_top.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/top/riscv_tcm_top.v"

`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/tcm/tcm_mem.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/tcm/tcm_mem_ram.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/tcm/tcm_mem_pmem.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/tcm/dport_axi.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/tcm/tcm_mem_rom.v"
`include "/home/altus/Cores-SweRV-EL2zybo/rtl/biriscv/tcm/dport_mux.v"

