`define VERILATOR

