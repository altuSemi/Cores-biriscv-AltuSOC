rom[0]=64'hba41819300002197;
rom[1]=64'hff81011300010117;
rom[2]=64'h1c40006f00010433;
rom[3]=64'h00112623ff010113;
rom[4]=64'h00f00313100012b7;
rom[5]=64'h00c120830062a823;
rom[6]=64'h0000806701010113;
rom[7]=64'h00112623ff010113;
rom[8]=64'h0142a303100012b7;
rom[9]=64'h0010039302058263;
rom[10]=64'h0010051300758663;
rom[11]=64'h00a343330240006f;
rom[12]=64'h0000051300628a23;
rom[13]=64'hfff545130140006f;
rom[14]=64'h00628a2300a37333;
rom[15]=64'h00c1208300000513;
rom[16]=64'h0000806701010113;
rom[17]=64'h00112623ff010113;
rom[18]=64'h00c1208300a58023;
rom[19]=64'h0000806701010113;
rom[20]=64'h00112623ff010113;
rom[21]=64'h100012b70004a303;
rom[22]=64'h0003a303005503b3;
rom[23]=64'h00c1208300030513;
rom[24]=64'h0000806701010113;
rom[25]=64'h00812e23fe010113;
rom[26]=64'hfea4262302010413;
rom[27]=64'hc0179073fec42783;
rom[28]=64'h01c1240300000013;
rom[29]=64'h0000806702010113;
rom[30]=64'h02112623fd010113;
rom[31]=64'h0301041302812423;
rom[32]=64'hfdc42783fca42e23;
rom[33]=64'hfe042623fef42423;
rom[34]=64'hc00027f30140006f;
rom[35]=64'hfe442783fef42223;
rom[36]=64'hfec42703fef42623;
rom[37]=64'hfef764e3fe842783;
rom[38]=64'hf95ff0ef00000513;
rom[39]=64'h02c1208300000013;
rom[40]=64'h0301011302812403;
rom[41]=64'hfe01011300008067;
rom[42]=64'h0201041300812e23;
rom[43]=64'hfec42703fea42623;
rom[44]=64'h04f70e6300800793;
rom[45]=64'h00800793fec42703;
rom[46]=64'hfec4270304e7cc63;
rom[47]=64'h02f70e6300400793;
rom[48]=64'h00400793fec42703;
rom[49]=64'hfec4270304e7c063;
rom[50]=64'h00f70a6300100793;
rom[51]=64'h00200793fec42703;
rom[52]=64'h0240006f00f70863;
rom[53]=64'h01c0006f00000793;
rom[54]=64'h0140006f00100793;
rom[55]=64'h00c0006f00200793;
rom[56]=64'h0040006f00300793;
rom[57]=64'h01c1240300078513;
rom[58]=64'h0000806702010113;
rom[59]=64'h02112e23fc010113;
rom[60]=64'h02912a2302812c23;
rom[61]=64'hfe04202304010413;
rom[62]=64'h36800793fe042623;
rom[63]=64'h0047a6830007a603;
rom[64]=64'h00c7a7830087a703;
rom[65]=64'hfcd42423fcc42223;
rom[66]=64'hfcf42823fce42623;
rom[67]=64'hfef4242300100793;
rom[68]=64'he7dff0ef01800513;
rom[69]=64'h0107979300050793;
rom[70]=64'h0017f7930107d793;
rom[71]=64'hfdc42783fcf42e23;
rom[72]=64'h0c80079300078863;
rom[73]=64'h0100006ffef42223;
rom[74]=64'h68078793009897b7;
rom[75]=64'hdbdff0effef42223;
rom[76]=64'he65ff0ef00000513;
rom[77]=64'hfe0426230dc0006f;
rom[78]=64'h014005130940006f;
rom[79]=64'h00050793e29ff0ef;
rom[80]=64'hfec42783fcf41d23;
rom[81]=64'hff04071300279793;
rom[82]=64'hfd47a78300f707b3;
rom[83]=64'h00078513fe842583;
rom[84]=64'h01400513d99ff0ef;
rom[85]=64'h00050793df9ff0ef;
rom[86]=64'hfda45703fcf41c23;
rom[87]=64'h00f747b3fd845783;
rom[88]=64'hfe842783fcf41b23;
rom[89]=64'hfd64178300479493;
rom[90]=64'he79ff0ef00078513;
rom[91]=64'h00f4873300050793;
rom[92]=64'h00878593100017b7;
rom[93]=64'hd9dff0ef00070513;
rom[94]=64'hdfdff0effe442503;
rom[95]=64'h00178793fec42783;
rom[96]=64'hfec42703fef42623;
rom[97]=64'hf6e7d4e300300793;
rom[98]=64'h00100793fe842703;
rom[99]=64'hfe04242300f71663;
rom[100]=64'h001007930240006f;
rom[101]=64'hfdc42783fef42423;
rom[102]=64'h100017b700078a63;
rom[103]=64'h0000051300978593;
rom[104]=64'hfe042783d49ff0ef;
rom[105]=64'h00000013f20782e3;
rom[106]=64'h03c1208300078513;
rom[107]=64'h0341248303812403;
rom[108]=64'h0000806704010113;
rom[109]=64'h0000000200000001;
rom[110]=64'h0000000800000004;
rom[111]=64'h0000000000000014;
rom[112]=64'h01017c0100527a03;
rom[113]=64'h0000000107020d1b;
rom[114]=64'h0000001c00000010;
rom[115]=64'h00000018fffffc68;
rom[116]=64'h0000000000000000
;
