`define VERILATOR
`define VIVADO

