`define VERILATOR
`define VIVADO
//`define AXI_HOST_IF

